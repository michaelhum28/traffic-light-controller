library verilog;
use verilog.vl_types.all;
entity Project_vlg_vec_tst is
end Project_vlg_vec_tst;
