library verilog;
use verilog.vl_types.all;
entity TXTEST_vlg_vec_tst is
end TXTEST_vlg_vec_tst;
