library verilog;
use verilog.vl_types.all;
entity COMP_TEST_vlg_check_tst is
    port(
        X               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end COMP_TEST_vlg_check_tst;
