library verilog;
use verilog.vl_types.all;
entity COUNTR_TEST_vlg_vec_tst is
end COUNTR_TEST_vlg_vec_tst;
