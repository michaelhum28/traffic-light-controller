library verilog;
use verilog.vl_types.all;
entity COUNTER_TEST_vlg_check_tst is
    port(
        \Out\           : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end COUNTER_TEST_vlg_check_tst;
