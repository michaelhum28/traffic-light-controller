library verilog;
use verilog.vl_types.all;
entity MUXTEST_vlg_vec_tst is
end MUXTEST_vlg_vec_tst;
