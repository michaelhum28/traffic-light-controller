library verilog;
use verilog.vl_types.all;
entity REGTEST_vlg_vec_tst is
end REGTEST_vlg_vec_tst;
