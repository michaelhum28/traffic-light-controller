library verilog;
use verilog.vl_types.all;
entity SUBXTEST_vlg_vec_tst is
end SUBXTEST_vlg_vec_tst;
