library verilog;
use verilog.vl_types.all;
entity TFF_TEST_vlg_vec_tst is
end TFF_TEST_vlg_vec_tst;
