library verilog;
use verilog.vl_types.all;
entity COMP_TEST_vlg_vec_tst is
end COMP_TEST_vlg_vec_tst;
