library verilog;
use verilog.vl_types.all;
entity FSMTEST_vlg_vec_tst is
end FSMTEST_vlg_vec_tst;
