library verilog;
use verilog.vl_types.all;
entity RXTEST_vlg_vec_tst is
end RXTEST_vlg_vec_tst;
