library verilog;
use verilog.vl_types.all;
entity MUXCT_TEST_vlg_vec_tst is
end MUXCT_TEST_vlg_vec_tst;
