library verilog;
use verilog.vl_types.all;
entity MUXTL_TEST_vlg_vec_tst is
end MUXTL_TEST_vlg_vec_tst;
